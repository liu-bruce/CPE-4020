'ifndef  Lab_3_libary.vh
'define Lab_3_libary.vh
module seven_segment_display_slot_6(light_segment_6, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_5(light_segment_5, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_4(light_segment_4, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_3(light_segment_3, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_2(light_segment_2, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_1(light_segment_1, input_a,input_b,input_c,input_d);
module seven_segment_display_slot_0(light_segment_0, input_a,input_b,input_c,input_d);
'endif
